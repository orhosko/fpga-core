
//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10.03 Education
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Mon Feb 17 17:27:46 2025

module Gowin_DPB (
    douta,
    doutb,
    clka,
    ocea,
    cea,
    reseta,
    wrea,
    clkb,
    oceb,
    ceb,
    resetb,
    wreb,
    ada,
    dina,
    adb,
    dinb
);

  output [7:0] douta;
  output [7:0] doutb;
  input clka;
  input ocea;
  input cea;
  input reseta;
  input wrea;
  input clkb;
  input oceb;
  input ceb;
  input resetb;
  input wreb;
  input [13:0] ada;
  input [7:0] dina;
  input [13:0] adb;
  input [7:0] dinb;

  wire [14:0] dpb_inst_0_douta_w;
  wire [14:0] dpb_inst_0_doutb_w;
  wire [14:0] dpb_inst_1_douta_w;
  wire [14:0] dpb_inst_1_doutb_w;
  wire [14:0] dpb_inst_2_douta_w;
  wire [14:0] dpb_inst_2_doutb_w;
  wire [14:0] dpb_inst_3_douta_w;
  wire [14:0] dpb_inst_3_doutb_w;
  wire [14:0] dpb_inst_4_douta_w;
  wire [14:0] dpb_inst_4_doutb_w;
  wire [14:0] dpb_inst_5_douta_w;
  wire [14:0] dpb_inst_5_doutb_w;
  wire [14:0] dpb_inst_6_douta_w;
  wire [14:0] dpb_inst_6_doutb_w;
  wire [14:0] dpb_inst_7_douta_w;
  wire [14:0] dpb_inst_7_doutb_w;
  wire gw_gnd;

  assign gw_gnd = 1'b0;

  DPB dpb_inst_0 (
      .DOA({dpb_inst_0_douta_w[14:0], douta[0]}),
      .DOB({dpb_inst_0_doutb_w[14:0], doutb[0]}),
      .CLKA(clka),
      .OCEA(ocea),
      .CEA(cea),
      .RESETA(reseta),
      .WREA(wrea),
      .CLKB(clkb),
      .OCEB(oceb),
      .CEB(ceb),
      .RESETB(resetb),
      .WREB(wreb),
      .BLKSELA({gw_gnd, gw_gnd, gw_gnd}),
      .BLKSELB({gw_gnd, gw_gnd, gw_gnd}),
      .ADA(ada[13:0]),
      .DIA({
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        dina[0]
      }),
      .ADB(adb[13:0]),
      .DIB({
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        dinb[0]
      })
  );

  defparam dpb_inst_0.READ_MODE0 = 1'b0; defparam dpb_inst_0.READ_MODE1 = 1'b0;
      defparam dpb_inst_0.WRITE_MODE0 = 2'b00; defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
      defparam dpb_inst_0.BIT_WIDTH_0 = 1; defparam dpb_inst_0.BIT_WIDTH_1 = 1;
      defparam dpb_inst_0.BLK_SEL_0 = 3'b000; defparam dpb_inst_0.BLK_SEL_1 = 3'b000;
      defparam dpb_inst_0.RESET_MODE = "SYNC";

  DPB dpb_inst_1 (
      .DOA({dpb_inst_1_douta_w[14:0], douta[1]}),
      .DOB({dpb_inst_1_doutb_w[14:0], doutb[1]}),
      .CLKA(clka),
      .OCEA(ocea),
      .CEA(cea),
      .RESETA(reseta),
      .WREA(wrea),
      .CLKB(clkb),
      .OCEB(oceb),
      .CEB(ceb),
      .RESETB(resetb),
      .WREB(wreb),
      .BLKSELA({gw_gnd, gw_gnd, gw_gnd}),
      .BLKSELB({gw_gnd, gw_gnd, gw_gnd}),
      .ADA(ada[13:0]),
      .DIA({
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        dina[1]
      }),
      .ADB(adb[13:0]),
      .DIB({
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        dinb[1]
      })
  );

  defparam dpb_inst_1.READ_MODE0 = 1'b0; defparam dpb_inst_1.READ_MODE1 = 1'b0;
      defparam dpb_inst_1.WRITE_MODE0 = 2'b00; defparam dpb_inst_1.WRITE_MODE1 = 2'b00;
      defparam dpb_inst_1.BIT_WIDTH_0 = 1; defparam dpb_inst_1.BIT_WIDTH_1 = 1;
      defparam dpb_inst_1.BLK_SEL_0 = 3'b000; defparam dpb_inst_1.BLK_SEL_1 = 3'b000;
      defparam dpb_inst_1.RESET_MODE = "SYNC";

  DPB dpb_inst_2 (
      .DOA({dpb_inst_2_douta_w[14:0], douta[2]}),
      .DOB({dpb_inst_2_doutb_w[14:0], doutb[2]}),
      .CLKA(clka),
      .OCEA(ocea),
      .CEA(cea),
      .RESETA(reseta),
      .WREA(wrea),
      .CLKB(clkb),
      .OCEB(oceb),
      .CEB(ceb),
      .RESETB(resetb),
      .WREB(wreb),
      .BLKSELA({gw_gnd, gw_gnd, gw_gnd}),
      .BLKSELB({gw_gnd, gw_gnd, gw_gnd}),
      .ADA(ada[13:0]),
      .DIA({
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        dina[2]
      }),
      .ADB(adb[13:0]),
      .DIB({
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        dinb[2]
      })
  );

  defparam dpb_inst_2.READ_MODE0 = 1'b0; defparam dpb_inst_2.READ_MODE1 = 1'b0;
      defparam dpb_inst_2.WRITE_MODE0 = 2'b00; defparam dpb_inst_2.WRITE_MODE1 = 2'b00;
      defparam dpb_inst_2.BIT_WIDTH_0 = 1; defparam dpb_inst_2.BIT_WIDTH_1 = 1;
      defparam dpb_inst_2.BLK_SEL_0 = 3'b000; defparam dpb_inst_2.BLK_SEL_1 = 3'b000;
      defparam dpb_inst_2.RESET_MODE = "SYNC";

  DPB dpb_inst_3 (
      .DOA({dpb_inst_3_douta_w[14:0], douta[3]}),
      .DOB({dpb_inst_3_doutb_w[14:0], doutb[3]}),
      .CLKA(clka),
      .OCEA(ocea),
      .CEA(cea),
      .RESETA(reseta),
      .WREA(wrea),
      .CLKB(clkb),
      .OCEB(oceb),
      .CEB(ceb),
      .RESETB(resetb),
      .WREB(wreb),
      .BLKSELA({gw_gnd, gw_gnd, gw_gnd}),
      .BLKSELB({gw_gnd, gw_gnd, gw_gnd}),
      .ADA(ada[13:0]),
      .DIA({
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        dina[3]
      }),
      .ADB(adb[13:0]),
      .DIB({
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        dinb[3]
      })
  );

  defparam dpb_inst_3.READ_MODE0 = 1'b0; defparam dpb_inst_3.READ_MODE1 = 1'b0;
      defparam dpb_inst_3.WRITE_MODE0 = 2'b00; defparam dpb_inst_3.WRITE_MODE1 = 2'b00;
      defparam dpb_inst_3.BIT_WIDTH_0 = 1; defparam dpb_inst_3.BIT_WIDTH_1 = 1;
      defparam dpb_inst_3.BLK_SEL_0 = 3'b000; defparam dpb_inst_3.BLK_SEL_1 = 3'b000;
      defparam dpb_inst_3.RESET_MODE = "SYNC";

  DPB dpb_inst_4 (
      .DOA({dpb_inst_4_douta_w[14:0], douta[4]}),
      .DOB({dpb_inst_4_doutb_w[14:0], doutb[4]}),
      .CLKA(clka),
      .OCEA(ocea),
      .CEA(cea),
      .RESETA(reseta),
      .WREA(wrea),
      .CLKB(clkb),
      .OCEB(oceb),
      .CEB(ceb),
      .RESETB(resetb),
      .WREB(wreb),
      .BLKSELA({gw_gnd, gw_gnd, gw_gnd}),
      .BLKSELB({gw_gnd, gw_gnd, gw_gnd}),
      .ADA(ada[13:0]),
      .DIA({
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        dina[4]
      }),
      .ADB(adb[13:0]),
      .DIB({
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        dinb[4]
      })
  );

  defparam dpb_inst_4.READ_MODE0 = 1'b0; defparam dpb_inst_4.READ_MODE1 = 1'b0;
      defparam dpb_inst_4.WRITE_MODE0 = 2'b00; defparam dpb_inst_4.WRITE_MODE1 = 2'b00;
      defparam dpb_inst_4.BIT_WIDTH_0 = 1; defparam dpb_inst_4.BIT_WIDTH_1 = 1;
      defparam dpb_inst_4.BLK_SEL_0 = 3'b000; defparam dpb_inst_4.BLK_SEL_1 = 3'b000;
      defparam dpb_inst_4.RESET_MODE = "SYNC";

  DPB dpb_inst_5 (
      .DOA({dpb_inst_5_douta_w[14:0], douta[5]}),
      .DOB({dpb_inst_5_doutb_w[14:0], doutb[5]}),
      .CLKA(clka),
      .OCEA(ocea),
      .CEA(cea),
      .RESETA(reseta),
      .WREA(wrea),
      .CLKB(clkb),
      .OCEB(oceb),
      .CEB(ceb),
      .RESETB(resetb),
      .WREB(wreb),
      .BLKSELA({gw_gnd, gw_gnd, gw_gnd}),
      .BLKSELB({gw_gnd, gw_gnd, gw_gnd}),
      .ADA(ada[13:0]),
      .DIA({
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        dina[5]
      }),
      .ADB(adb[13:0]),
      .DIB({
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        dinb[5]
      })
  );

  defparam dpb_inst_5.READ_MODE0 = 1'b0; defparam dpb_inst_5.READ_MODE1 = 1'b0;
      defparam dpb_inst_5.WRITE_MODE0 = 2'b00; defparam dpb_inst_5.WRITE_MODE1 = 2'b00;
      defparam dpb_inst_5.BIT_WIDTH_0 = 1; defparam dpb_inst_5.BIT_WIDTH_1 = 1;
      defparam dpb_inst_5.BLK_SEL_0 = 3'b000; defparam dpb_inst_5.BLK_SEL_1 = 3'b000;
      defparam dpb_inst_5.RESET_MODE = "SYNC";

  DPB dpb_inst_6 (
      .DOA({dpb_inst_6_douta_w[14:0], douta[6]}),
      .DOB({dpb_inst_6_doutb_w[14:0], doutb[6]}),
      .CLKA(clka),
      .OCEA(ocea),
      .CEA(cea),
      .RESETA(reseta),
      .WREA(wrea),
      .CLKB(clkb),
      .OCEB(oceb),
      .CEB(ceb),
      .RESETB(resetb),
      .WREB(wreb),
      .BLKSELA({gw_gnd, gw_gnd, gw_gnd}),
      .BLKSELB({gw_gnd, gw_gnd, gw_gnd}),
      .ADA(ada[13:0]),
      .DIA({
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        dina[6]
      }),
      .ADB(adb[13:0]),
      .DIB({
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        dinb[6]
      })
  );

  defparam dpb_inst_6.READ_MODE0 = 1'b0; defparam dpb_inst_6.READ_MODE1 = 1'b0;
      defparam dpb_inst_6.WRITE_MODE0 = 2'b00; defparam dpb_inst_6.WRITE_MODE1 = 2'b00;
      defparam dpb_inst_6.BIT_WIDTH_0 = 1; defparam dpb_inst_6.BIT_WIDTH_1 = 1;
      defparam dpb_inst_6.BLK_SEL_0 = 3'b000; defparam dpb_inst_6.BLK_SEL_1 = 3'b000;
      defparam dpb_inst_6.RESET_MODE = "SYNC";

  DPB dpb_inst_7 (
      .DOA({dpb_inst_7_douta_w[14:0], douta[7]}),
      .DOB({dpb_inst_7_doutb_w[14:0], doutb[7]}),
      .CLKA(clka),
      .OCEA(ocea),
      .CEA(cea),
      .RESETA(reseta),
      .WREA(wrea),
      .CLKB(clkb),
      .OCEB(oceb),
      .CEB(ceb),
      .RESETB(resetb),
      .WREB(wreb),
      .BLKSELA({gw_gnd, gw_gnd, gw_gnd}),
      .BLKSELB({gw_gnd, gw_gnd, gw_gnd}),
      .ADA(ada[13:0]),
      .DIA({
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        dina[7]
      }),
      .ADB(adb[13:0]),
      .DIB({
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        gw_gnd,
        dinb[7]
      })
  );

  defparam dpb_inst_7.READ_MODE0 = 1'b0; defparam dpb_inst_7.READ_MODE1 = 1'b0;
      defparam dpb_inst_7.WRITE_MODE0 = 2'b00; defparam dpb_inst_7.WRITE_MODE1 = 2'b00;
      defparam dpb_inst_7.BIT_WIDTH_0 = 1; defparam dpb_inst_7.BIT_WIDTH_1 = 1;
      defparam dpb_inst_7.BLK_SEL_0 = 3'b000; defparam dpb_inst_7.BLK_SEL_1 = 3'b000;
      defparam dpb_inst_7.RESET_MODE = "SYNC";

endmodule  //Gowin_DPB

